`timescale 1ns/1ns

module tb_top_scope;

    //==========================================================================
    // 1. �źŶ���
    //==========================================================================
    reg             sys_clk;
    reg             sys_rst_n;
    reg     [7:0]   ad_data;    // ģ��ADC����
    reg             key_start;  // ����1
    reg             key_mode;   // ����2

    wire            ad_clk;     // �����ADC��ʱ��
    wire    [5:0]   sel;        // �����λѡ
    wire    [7:0]   seg;        // ����ܶ�ѡ

    // ���������������������ǲ�
    reg             dir;        // 0: ��������, 1: ��������
    
    //==========================================================================
    // 2. ģ��ʵ���� (DUT - Device Under Test)
    //==========================================================================
    top_scope uut (
        .sys_clk    (sys_clk),
        .sys_rst_n  (sys_rst_n),
        .ad_data    (ad_data),
        .key_start  (key_start),
        .key_mode   (key_mode),
        .ad_clk     (ad_clk),
        .sel        (sel),
        .seg        (seg)
    );

    //==========================================================================
    // 3. ������д (Ϊ���÷����ܵÿ죬�����޸���Щ������)
    //==========================================================================
    // ע�⣺�����·����������ģ��ʵ��������һ��
    
    // ���̰�������ʱ�� (ԭ20ms -> ��Ϊ4��ʱ������)
    defparam uut.key_start_inst.CNT_MAX = 20'd4;
    defparam uut.key_mode_inst.CNT_MAX  = 20'd4;
    
    // ����ADCУ׼ʱ�� (ԭ1024�� -> ��Ϊ64��)
    defparam uut.adc_inst.CNT_DATA_MAX  = 11'd64;

    // ���̷�ֵ���ˢ��ʱ�� (ԭ0.3�� -> ��Ϊ2000��ʱ��)
    defparam uut.CNT_PEAK_MAX           = 25'd2000;
    
    // ����Ƶ�ʼ�բ��ʱ�� (ԭ1�� -> ��Ϊ4000��ʱ��)
    defparam uut.freq_meter_inst.CNT_1S_MAX = 26'd4000;

    //==========================================================================
    // 4. ʱ������ (50MHz)
    //==========================================================================
    initial begin
        sys_clk = 0;
        forever #10 sys_clk = ~sys_clk; // 20ns����
    end

    //==========================================================================
    // 5. ���ݷ��������������ǲ� (ģ��仯�ĵ�ѹ)
    //==========================================================================
    // �߼����� ad_clk ���½��ظ������ݣ�ģ�� ADC оƬ��Ϊ
    always @(negedge ad_clk or negedge sys_rst_n) begin
        if(!sys_rst_n) begin
            ad_data <= 8'd128; // ��λ�����ֵ
            dir     <= 0;
        end 
        else if (uut.adc_inst.median_en == 1'b0) begin
            // У׼�ڼ䣬�����ȶ�����ֵ���� (ģ��0V)
            ad_data <= 8'd128;
        end
        else begin
            // У׼��ɺ��������ǲ� (0 -> 255 -> 0)
            if(dir == 0) begin
                if(ad_data >= 8'd254) dir <= 1;
                else ad_data <= ad_data + 1;
            end else begin
                if(ad_data <= 8'd1)   dir <= 0;
                else ad_data <= ad_data - 1;
            end
        end
    end

    //==========================================================================
    // 6. �������� (���߾���)
    //==========================================================================
    initial begin
        // --- ��ʼ�� ---
        sys_rst_n = 0;
        key_start = 1; // ����δ����(�ߵ�ƽ)
        key_mode  = 1;
        $display("--------------------------------------------------");
        $display("Simulation Start: System Reset");
        $display("--------------------------------------------------");

        // --- �ͷŸ�λ ---
        #200;
        sys_rst_n = 1;
        
        // --- �ȴ� ADC �Զ�У׼��� ---
        $display("Status: Waiting for ADC Auto-Calibration...");
        wait(uut.adc_inst.median_en == 1'b1);
        $display("Status: ADC Calibration Done! Zero-point set at %d", uut.adc_inst.data_median);
        
        // --- ��ʱ��Ȼ�в������룬��ϵͳ����PAUSE״̬�������Ӧ��ʾ0�򲻸��� ---
        #1000;

        // --- ����1�����¿�ʼ�� (Start) ---
        $display("Action: Pressing START Key...");
        key_start = 0; #100; // ����
        key_start = 1; #100; // �ͷ�
        
        // --- ����һ��ʱ�䣬�۲��ֵ���� ---
        // ���������ǲ�(0~255)����ֵӦ�ñ���׽����ʾ
        $display("Status: System Running... Monitoring Peak Voltage...");
        #60000; 

        // --- ����2������ģʽ�� (Mode Switch) ---
        $display("Action: Pressing MODE Key (Switch to Frequency)...");
        key_mode = 0; #100;
        key_mode = 1; #100;

        // --- ����һ��ʱ�䣬�۲�Ƶ����ʾ ---
        $display("Status: Mode Switched. Measuring Frequency...");
        #60000;

        // --- �������� ---
        $display("--------------------------------------------------");
        $display("Simulation Finished.");
        $display("--------------------------------------------------");
        $stop; 
    end

    //==========================================================================
    // 7. ʵʱ��ش�ӡ (Debug helper)
    //==========================================================================
    // ÿ�� 5000ns ��ӡһ�ιؼ�״̬����ֹ�㶢�ſհ���Ļ����
    always begin
        #5000;
        if($time > 200) begin
            $display("Time: %t | State: %s | ADC_Raw: %d | Volt_Inst: %d mV | Disp_Peak: %d mV | Freq: %d Hz", 
                     $time, 
                     (uut.run_state ? "RUN " : "STOP"), 
                     ad_data, 
                     uut.volt_inst, 
                     uut.volt_display,
                     uut.freq_val);
        end
    end

endmodule